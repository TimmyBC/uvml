class eg_hs_seq extends uvml_sequence;
    
//    static function eg_hs_seq create(string name);
//        eg_hs_seq seq = new(name);
//        return seq;
//    endfunction
    
    function new(string name);
        super.new(name);
    endfunction
    
endclass : eg_hs_seq
