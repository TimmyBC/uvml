package uvml_stream_pkg;
    import uvml_pkg::*;
    import uvml_hs_pkg::*;
    `include "uvml_macros.svh"
    
    `include "uvml_stream_drive_pattern.svh"
    `include "uvml_stream_if_api.svh"
    `include "uvml_stream_seq_item.svh"
    `include "uvml_stream_packer.svh"
    `include "uvml_stream_monitor.svh"
    `include "uvml_stream_driver.svh"
    `include "uvml_stream_agent.svh"
endpackage
