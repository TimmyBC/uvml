package uvml_hs_pkg;
	import uvml_pkg::*;
	`include "uvml_macros.svh"
    
    `include "uvml_hs_drive_pattern.svh"
    `include "uvml_hs_if_api.svh"
	`include "uvml_hs_seq_item.svh"
    `include "uvml_hs_packer.svh"
//    typedef uvml_api_sequence#(T) uvml_hs_api_sequence#(T);
	`include "uvml_hs_monitor.svh"
	`include "uvml_hs_driver.svh"
	`include "uvml_hs_agent.svh"
endpackage
