class uvml_monitor extends uvml_component;

	function new(string name, uvml_component parent);
		super.new(name, parent);
		
	endfunction

endclass : uvml_monitor
